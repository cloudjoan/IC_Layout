* SPICE NETLIST
***************************************

.SUBCKT CLKINVX1
** N=4 EP=0 IP=0 FDC=2
M0 3 4 2 2 nmos1v L=1e-07 W=4.3e-07 $X=235 $Y=325 $D=5
M1 3 4 1 1 pmos1v L=1e-07 W=6.5e-07 $X=235 $Y=1230 $D=6
.ENDS
***************************************

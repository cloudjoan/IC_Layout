* SPICE NETLIST
***************************************

.SUBCKT INVX16 VDD VSS Y A
** N=4 EP=4 IP=0 FDC=32
M0 Y A VSS VSS nmos1v L=1e-07 W=4.3e-07 $X=280 $Y=1825 $D=5
M1 VSS A Y VSS nmos1v L=1e-07 W=4.3e-07 $X=720 $Y=1825 $D=5
M2 Y A VSS VSS nmos1v L=1e-07 W=4.3e-07 $X=1155 $Y=1825 $D=5
M3 VSS A Y VSS nmos1v L=1e-07 W=4.3e-07 $X=1600 $Y=1825 $D=5
M4 Y A VSS VSS nmos1v L=1e-07 W=4.3e-07 $X=2040 $Y=1825 $D=5
M5 VSS A Y VSS nmos1v L=1e-07 W=4.3e-07 $X=2475 $Y=1825 $D=5
M6 Y A VSS VSS nmos1v L=1e-07 W=4.3e-07 $X=2920 $Y=1825 $D=5
M7 VSS A Y VSS nmos1v L=1e-07 W=4.3e-07 $X=3350 $Y=1825 $D=5
M8 Y A VSS VSS nmos1v L=1e-07 W=4.3e-07 $X=3780 $Y=1825 $D=5
M9 VSS A Y VSS nmos1v L=1e-07 W=4.3e-07 $X=4220 $Y=1825 $D=5
M10 Y A VSS VSS nmos1v L=1e-07 W=4.3e-07 $X=4655 $Y=1825 $D=5
M11 VSS A Y VSS nmos1v L=1e-07 W=4.3e-07 $X=5100 $Y=1825 $D=5
M12 Y A VSS VSS nmos1v L=1e-07 W=4.3e-07 $X=5540 $Y=1825 $D=5
M13 VSS A Y VSS nmos1v L=1e-07 W=4.3e-07 $X=5975 $Y=1825 $D=5
M14 Y A VSS VSS nmos1v L=1e-07 W=4.3e-07 $X=6420 $Y=1825 $D=5
M15 VSS A Y VSS nmos1v L=1e-07 W=4.3e-07 $X=6850 $Y=1825 $D=5
M16 Y A VDD VDD pmos1v L=1e-07 W=6.5e-07 $X=280 $Y=2765 $D=6
M17 VDD A Y VDD pmos1v L=1e-07 W=6.5e-07 $X=720 $Y=2765 $D=6
M18 Y A VDD VDD pmos1v L=1e-07 W=6.5e-07 $X=1150 $Y=2765 $D=6
M19 VDD A Y VDD pmos1v L=1e-07 W=6.5e-07 $X=1595 $Y=2765 $D=6
M20 Y A VDD VDD pmos1v L=1e-07 W=6.5e-07 $X=2035 $Y=2765 $D=6
M21 VDD A Y VDD pmos1v L=1e-07 W=6.5e-07 $X=2465 $Y=2765 $D=6
M22 Y A VDD VDD pmos1v L=1e-07 W=6.5e-07 $X=2915 $Y=2765 $D=6
M23 VDD A Y VDD pmos1v L=1e-07 W=6.5e-07 $X=3345 $Y=2765 $D=6
M24 Y A VDD VDD pmos1v L=1e-07 W=6.5e-07 $X=3780 $Y=2765 $D=6
M25 VDD A Y VDD pmos1v L=1e-07 W=6.5e-07 $X=4220 $Y=2765 $D=6
M26 Y A VDD VDD pmos1v L=1e-07 W=6.5e-07 $X=4650 $Y=2765 $D=6
M27 VDD A Y VDD pmos1v L=1e-07 W=6.5e-07 $X=5095 $Y=2765 $D=6
M28 Y A VDD VDD pmos1v L=1e-07 W=6.5e-07 $X=5535 $Y=2765 $D=6
M29 VDD A Y VDD pmos1v L=1e-07 W=6.5e-07 $X=5965 $Y=2765 $D=6
M30 Y A VDD VDD pmos1v L=1e-07 W=6.5e-07 $X=6415 $Y=2765 $D=6
M31 VDD A Y VDD pmos1v L=1e-07 W=6.5e-07 $X=6845 $Y=2765 $D=6
.ENDS
***************************************
